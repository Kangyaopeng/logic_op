`ifndef TB_CLK_DIVIDER__SV
`define TB_CLK_DIVIDER__SV
module tb_clk_div #(parameter WIDTH = 3, parameter DIV_NUM = 6)
              (
		            input  clk,
		            input  rst_n,
		            output o_clk
		          );

endmodule
`endif
