`ifndef LOGIC_OP_DEFINE__SV
`define LOGIC_OP_DEFINE__SV

//  `define ABC abc
//  `define BCD
  //`ifdef RUN_LOGIC_OP
    `define MERGE_ITF_NAME(prename, name) prename``name
    `define LOGIC_OP_PATH logic_op_tb_top.u_logic_op
    `define REG_UPD_ADDR 32'h4000_0004

    //-----------------------------------------------------------
    //-----------------------------------------------------------

    //Sub Env Define
  //`endif

`endif
