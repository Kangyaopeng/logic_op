`ifndef OP_IN_SEQ_PACKAGE__SV
`define OP_IN_SEQ_PACKAGE__SV
package op_in_seq_pkg;
  import uvm_pkg::*;

  `include "op_in_seq_lib.svh"

endpackage
`endif
