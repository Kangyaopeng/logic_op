package logic_reg_model_pkg;
  import uvm_pkg::*;
  //sub-reg_model pkg
  `include "logic_reg_field.svh"
  `include "logic_reg_model.svh"
endpackage
