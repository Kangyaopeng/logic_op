`ifndef OP_OUT_SEQ_PACKAGE__SV
`define OP_OUT_SEQ_PACKAGE__SV
package op_out_seq_pkg;
  import uvm_pkg::*;

  `include "op_out_seq_lib.svh"

endpackage
`endif
