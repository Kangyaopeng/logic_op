`ifndef OP_OUT_AGENT_PACKAGE__SV
`define OP_OUT_AGENT_PACKAGE__SV
package op_out_agent_pkg;

import uvm_pkg::*;

`include "op_out_agent_config.svh"
`include "op_out_seq_item.svh"
`include "op_out_driver.svh"
`include "op_out_monitor.svh"
`include "op_out_sequencer.svh"
`include "op_out_agent.svh"

//adapter here

`include "op_out_seq_lib.svh"

endpackage

`include "op_out_if.sv"

  

`endif
